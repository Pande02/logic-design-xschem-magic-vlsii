magic
tech sky130A
magscale 1 2
timestamp 1729065313
<< metal1 >>
rect 146 2312 606 2313
rect 146 2272 1030 2312
rect 146 2200 188 2272
rect 565 2271 1030 2272
rect 565 2192 606 2271
rect 989 2188 1030 2271
rect 126 1838 204 1844
rect 126 1786 136 1838
rect 190 1786 204 1838
rect 1128 1838 1220 1846
rect 286 1798 661 1828
rect 710 1800 1038 1828
rect 126 1780 204 1786
rect 1128 1786 1144 1838
rect 1204 1786 1220 1838
rect 1128 1776 1220 1786
rect 140 1354 184 1452
rect 558 1354 604 1428
rect 986 1354 1030 1446
rect 140 1310 1030 1354
<< via1 >>
rect 136 1786 190 1838
rect 1144 1786 1204 1838
<< metal2 >>
rect 130 1840 200 1844
rect 1136 1840 1214 1844
rect 130 1838 1214 1840
rect 130 1786 136 1838
rect 190 1786 1144 1838
rect 1204 1786 1214 1838
rect 130 1780 200 1786
rect 1136 1780 1214 1786
use modul_inv  x1 ~/MSIB/inverter
timestamp 1729064850
transform 1 0 53 0 1 1306
box -54 -53 369 1074
use modul_inv  x2
timestamp 1729064850
transform 1 0 474 0 1 1305
box -54 -53 369 1074
use modul_inv  x3
timestamp 1729064850
transform 1 0 896 0 1 1305
box -54 -53 369 1074
<< labels >>
flabel metal1 586 1330 586 1330 0 FreeSans 160 0 0 0 GND
port 2 nsew
flabel metal1 590 2288 590 2288 0 FreeSans 160 0 0 0 VDD
port 1 nsew
flabel metal2 638 1812 638 1812 0 FreeSans 160 0 0 0 OUT
port 3 nsew
<< end >>
